Vsource vin 0 DC 12
R1 vin vout 1k
R2 vout 0 470

.control
tran .5s 1s
.endc
.end
