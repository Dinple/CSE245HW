* netlist
V1 n1 0 SIN(0 1 6Hz)
C1 n2 0 1
R1 n2 n1 1
L1 0 n2 1
.END